TLM Communications
Blocking and Non-blocking ports
PUT port
GET port
Transport port
Analysis Port
TLM FIFO


