//* 1. Configuring TB env
//* 2. System Reset
//* 3. Applying Stimulus to DUT
//* 4. Comparing Response with Golden Data
//* 5. Generating Report

