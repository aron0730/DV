semaphore 	[identifier_name];

