// The super keyword is used from within a sub-class to refer to properties and methods of the base class

// Example
