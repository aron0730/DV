`timescale 1ns/1ps

module tb();
    
endmodule