module tb_and;
    

endmodule