Sequences
Sending Transactions to Driver
Multiple Sequences in Parallel
Arbitration Mechanism
Lock-Unlock Method
Grab-Ungrab Method