module dut(
    input [3:0] a, b,
    output [3:0] y
);


endmodule