// Step1: Callback Class
class MyCallback;
    virtual function void callback_function();
        // Default implementation (optional)
    endfunction
endclass