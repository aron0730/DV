// Syntax
/*
function int $cast (targ_var, source_exp);

task $cast (targ_var, source_exp);
*/

// Example
