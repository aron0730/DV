module fifo (
    input wreq, rreq,
    input clk,
    input rst,
    input [7:0] wdata,
    output [7:0] rdata,
    output full, empty;
);


endmodule