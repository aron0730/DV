module tb;

    initial
        $display("Hello world ! ");
endmodule