// Syntax
[default] clocking [identifier_name] @ [event_or_identifier]
    default input #[delay_or_edge] output #[delay_or_edge]
    [list of signals]
endclocking

