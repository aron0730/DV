Sequencer -> Driver : Special TLM Port : SEQ_ITEM_PORT

Monitor -> Scoreboard : TLP PORT : UVM_ANALYSIS PORT